module ALU (operand1, operand2, opSel, result,zero );
	parameter data_width = 32;
	parameter sel_width = 4;
	//input for alu
	input [data_width - 1 : 0] operand1, operand2;
	//selector to select operation
	input [sel_width - 1 :0] opSel;
	//output
	output reg [data_width - 1 : 0] result;
	output reg zero;
	
	parameter   	_ADD  = 4'b0000,
 			_SUB  = 4'b0001,
			_AND  = 4'b0010, 
			_OR   = 4'b0011,
			_NOR  = 4'b0100,
			_XOR  = 4'b0101,     
			_SLT  = 4'b0110,
			_SLL  = 4'b0111,
			_SRL  = 4'b1000,
			_SGT  = 4'b1001;

	always @ (*) begin
		case(opSel)
			_ADD: result = operand1 + operand2;
			_SUB: result = operand1 - operand2;
			_AND: result = operand1 & operand2;
			_OR: result = operand1 | operand2;
			_NOR: result = ~(operand1 | operand2);
			_XOR: result = operand1 ^ operand2;
			_SLT: result = (operand1 < operand2) ? 1 : 0; 
			_SLL: result = (operand1 << operand2[10:6]);
			_SRL: result = (operand1 >> operand2[10:6]);
			_SGT: result = (operand1 > operand2) ? 1 : 0;
			default : result = 32'b0 ;
		endcase
	end
	
	always @ (*) begin 
		
		zero = (result == 'b0);
	
	end

endmodule