module ANDGate(in1, in2, out);
	//input
	input in1, in2;
	//output
	output out;
	
	assign out = in1 & in2;
	
endmodule
